/*
*Author : Revanth Sai Nandamuri
*GitHUB : https://github.com/RevanthNandamuri1341b0
*Date of update : 29 July 2021
*Time of update : 15:29
*Project name : Router 4x4 Verification
*Domain : UVM
*Description : Sequence [SA1 -> Rest all OP ports]
File Name : sa1_sequence.sv
*File ID : 670073
*Modified by : #your name#
*/

class sa1_sequence extends uvm_sequence#(packet);
    int unsigned item_count;
    `uvm_object_utils(sa1_sequence);

    function new(string name = "sa1_sequence");
        super.new(name);
        set_automatic_phase_objection(1);
    endfunction: new

    extern virtual task pre_start();
    extern virtual task body();
    
endclass: sa1_sequence

task sa1_sequence::pre_start();
    if(!uvm_config_db #(int)::get(get_sequencer(),"","item_count",item_count))
    begin
        `uvm_warning(get_full_name(),"item_count is not set in sa1_sequencer");
        item_count=10;
    end
endtask: pre_start

task sa1_sequence::body();
    bit[31:0]count;
    REQ ref_pkt;
    ref_pkt=packet::type_id::create("ref_pkt",,get_full_name());
    repeat(item_count)
    begin
        `uvm_create(req);
        assert(ref_pkt.randomize() with {sa==1;});
        req.copy(ref_pkt);
        req.mode=STIMULUS;
        start_item(req);
        finish_item(req);
        count++;
        `uvm_info("SEQ",$sformatf("MASTER SEQUENCE : Transaction %0d DONE ",count ), UVM_MEDIUM);
    end
endtask: body
