/*
*Author : Revanth Sai Nandamuri
*GitHUB : https://github.com/RevanthNandamuri1341b0
*Date of update : 29 July 2021
*Time of update : 15:50
*Project name : Router 4x4 Verification
*Domain : UVM
*Description : Sequencer file to send sequence of stimulus
File Name : sequencer.sv
*File ID : 398975
*Modified by : #your name#
*/

typedef uvm_sequencer #(packet) sequencer;